module InstructionMemory(input [7:0] pc, output wire [15:0] instruction,output wire[15:0] next_instruction );  
     reg [15:0] rom[255:0];  
     initial  begin  
          rom[8'd0]  = 16'b0001_0000_0001_0010;  
          rom[8'd1]  = 16'b0001_0000_0001_0011;  
          rom[8'd2]  = 16'b0001_0000_1011_0100;  
          rom[8'd3]  = 16'b1000_0010_0011_0010;  
          rom[8'd4]  = 16'b0110_0010_0100_0110;  
          rom[8'd5]  = 16'b0000_0000_0000_0111; 
          rom[8'd6]  = 16'b0101_0000_0000_0011;  
          rom[8'd7]  = 16'b0000000000000000;  
          rom[8'd8]  = 16'b0000000000000000;  
          rom[8'd9]  = 16'b0000000000000000;  
          rom[8'd10] = 16'b0000000000000000;  
          rom[8'd11] = 16'b0000000000000000;  
          rom[8'd12] = 16'b0000000000000000;  
          rom[8'd13] = 16'b0000000000000000;  
          rom[8'd14] = 16'b0000000000000000;  
          rom[8'd15] = 16'b0000000000000000; 
          rom[8'd16] = 16'b0000000000000000; 
          rom[8'd17] = 16'b0000000000000000;   
          rom[8'd18] = 16'b0000000000000000;  
          rom[8'd19] = 16'b0000000000000000;  
          rom[8'd20] = 16'b0000000000000000;  
          rom[8'd21] = 16'b0000000000000000;  
          rom[8'd22] = 16'b0000000000000000;  
          rom[8'd23] = 16'b0000000000000000;  
          rom[8'd24] = 16'b0000000000000000;  
          rom[8'd25] = 16'b0000000000000000;  
          rom[8'd26] = 16'b0000000000000000;  
          rom[8'd27] = 16'b0000000000000000;  
          rom[8'd28] = 16'b0000000000000000;  
          rom[8'd29] = 16'b0000000000000000;  
          rom[8'd30] = 16'b0000000000000000;  
          rom[8'd31] = 16'b0000000000000000;  
          rom[8'd32] = 16'b0000000000000000;  
     end  
     assign instruction = (pc < 32 )? rom[pc]: 16'd0;  
     assign next_instruction = (pc < 31 )? rom[pc+1]: 16'd0;  
 endmodule   